library ieee;
use ieee.std_logic_1164.all;

entity can_generator is
  port (channel_0 : out std_ulogic);
end entity can_generator;

architecture tb of can_generator is
begin
  stimuli_proc : process
  begin
channel_0 <= '1';
wait for 46720 ns;
channel_0 <= '0';
wait for 10020 ns;
channel_0 <= '1';
wait for 1980 ns;
channel_0 <= '0';
wait for 10020 ns;
channel_0 <= '1';
wait for 1980 ns;
channel_0 <= '0';
wait for 2020 ns;
channel_0 <= '1';
wait for 1980 ns;
channel_0 <= '0';
wait for 6020 ns;
channel_0 <= '1';
wait for 1980 ns;
channel_0 <= '0';
wait for 10020 ns;
channel_0 <= '1';
wait for 1980 ns;
channel_0 <= '0';
wait for 10020 ns;
channel_0 <= '1';
wait for 3980 ns;
channel_0 <= '0';
wait for 10020 ns;
channel_0 <= '1';
wait for 1980 ns;
channel_0 <= '0';
wait for 4020 ns;
channel_0 <= '1';
wait for 1980 ns;
channel_0 <= '0';
wait for 6020 ns;
channel_0 <= '1';
wait for 1980 ns;
channel_0 <= '0';
wait for 2020 ns;
channel_0 <= '1';
wait for 1980 ns;
channel_0 <= '0';
wait for 2020 ns;
channel_0 <= '1';
wait for 1980 ns;
channel_0 <= '0';
wait for 10020 ns;
channel_0 <= '1';
wait for 1980 ns;
channel_0 <= '0';
wait for 10020 ns;
channel_0 <= '1';
wait for 1980 ns;
channel_0 <= '0';
wait for 10020 ns;
channel_0 <= '1';
wait for 1980 ns;
channel_0 <= '0';
wait for 10020 ns;
channel_0 <= '1';
wait for 1980 ns;
channel_0 <= '0';
wait for 10020 ns;
channel_0 <= '1';
wait for 1980 ns;
channel_0 <= '0';
wait for 10020 ns;
channel_0 <= '1';
wait for 1980 ns;
channel_0 <= '0';
wait for 10020 ns;
channel_0 <= '1';
wait for 1979 ns;
channel_0 <= '0';
wait for 10021 ns;
channel_0 <= '1';
wait for 1980 ns;
channel_0 <= '0';
wait for 2020 ns;
channel_0 <= '1';
wait for 3980 ns;
channel_0 <= '0';
wait for 6020 ns;
channel_0 <= '1';
wait for 1980 ns;
channel_0 <= '0';
wait for 2020 ns;
channel_0 <= '1';
wait for 3980 ns;
channel_0 <= '0';
wait for 2020 ns;
channel_0 <= '1';
wait for 10000 ns;
    wait;
  end process;
end architecture;
