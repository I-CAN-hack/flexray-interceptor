library ieee;
use ieee.std_logic_1164.all;

entity flexray_generator is
  port (channel_0 : out std_ulogic);
end entity flexray_generator;

architecture tb of flexray_generator is
begin
  stimuli_proc : process
  begin

wait for 10000 ns;
channel_0 <= '1';
wait for 10000 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 140 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8770 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9120 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9440 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9020 ns;
channel_0 <= '0';
wait for 940 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8680 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 140 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8750 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 113570 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 8870 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 166020 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9320 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9300 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 61330 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9220 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9270 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61190 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9050 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61470 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61660 ns;
channel_0 <= '0';
wait for 739 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 311 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 399 ns;
channel_0 <= '0';
wait for 401 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 8790 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 399 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 389 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 165929 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 799 ns;
channel_0 <= '1';
wait for 61601 ns;
channel_0 <= '0';
wait for 739 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 501 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 401 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 165441 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 209 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 211 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 289 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 311 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 491 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 191 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 591 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 311 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 309 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 409 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 309 ns;
channel_0 <= '0';
wait for 191 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 191 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 211 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 391 ns;
channel_0 <= '1';
wait for 9230 ns;
channel_0 <= '0';
wait for 939 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 501 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 401 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 599 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8960 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 599 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 599 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 799 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 701 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 401 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 108450 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 1601 ns;
channel_0 <= '1';
wait for 18270 ns;
channel_0 <= '0';
wait for 749 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 399 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 399 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 599 ns;
channel_0 <= '1';
wait for 1000000 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9440 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 9130 ns;
channel_0 <= '0';
wait for 940 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 120 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8570 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8750 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 9100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 113980 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 8790 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 166010 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9410 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9330 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 61210 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9270 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 610 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 9240 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9270 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61140 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9050 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61490 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 61760 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 8670 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 165950 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 61660 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 165360 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 45100 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 7600 ns;
channel_0 <= '1';
wait for 63370 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 18350 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1600 ns;
channel_0 <= '1';
wait for 342000 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 3600 ns;
channel_0 <= '1';
wait for 1000000 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9470 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 8990 ns;
channel_0 <= '0';
wait for 940 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 120 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8670 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9080 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 113880 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 8890 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 166030 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 290 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 610 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9300 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9320 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 61350 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9150 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9270 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61260 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9050 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 61460 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 710 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9220 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 1000 ns;
channel_0 <= '1';
wait for 61690 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 8790 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 165920 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61600 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 165460 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8780 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 560 ns;
channel_0 <= '1';
wait for 9580 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 90260 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 18460 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1600 ns;
channel_0 <= '1';
wait for 18230 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 99460 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1600 ns;
channel_0 <= '1';
wait for 45010 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 3590 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 1000000 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 420 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 220 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 9460 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 940 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8570 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9080 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 113630 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 8810 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 166020 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9380 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 9340 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61250 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9200 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 610 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 9270 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61230 ns;
channel_0 <= '0';
wait for 960 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9040 ns;
channel_0 <= '0';
wait for 960 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 61420 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9230 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 61780 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 8690 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 165910 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61680 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 165380 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8780 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 570 ns;
channel_0 <= '1';
wait for 140 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 98880 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 120 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 120 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 140 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 18230 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1600 ns;
channel_0 <= '1';
wait for 108360 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 6570 ns;
channel_0 <= '1';
wait for 9370 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 610 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 2600 ns;
channel_0 <= '1';
wait for 225070 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 3570 ns;
channel_0 <= '1';
wait for 1000000 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8790 ns;
channel_0 <= '0';
wait for 880 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 9100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 140 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 9130 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9000 ns;
channel_0 <= '0';
wait for 940 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 120 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8680 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9080 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8780 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 113880 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 8890 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 166060 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9280 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9310 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61350 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 9210 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 9270 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61210 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9040 ns;
channel_0 <= '0';
wait for 960 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61440 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9230 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 61690 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 8790 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 165900 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61620 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 165460 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9390 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 610 ns;
channel_0 <= '1';
wait for 36410 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 7590 ns;
channel_0 <= '1';
wait for 63430 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 580 ns;
channel_0 <= '1';
wait for 18320 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1600 ns;
channel_0 <= '1';
wait for 18230 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 710 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 390 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 90120 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 9560 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1600 ns;
channel_0 <= '1';
wait for 1000000 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 140 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8780 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9450 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9120 ns;
channel_0 <= '0';
wait for 940 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 810 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8570 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 9080 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 113640 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 8810 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 166080 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9340 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9310 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61260 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9270 ns;
channel_0 <= '0';
wait for 720 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9240 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9280 ns;
channel_0 <= '0';
wait for 720 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61160 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9050 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61440 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9230 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 61780 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 8710 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 165890 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61710 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 165380 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9650 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 18280 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 81240 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 18340 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1600 ns;
channel_0 <= '1';
wait for 108020 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 920 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 570 ns;
channel_0 <= '1';
wait for 234220 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 3600 ns;
channel_0 <= '1';
wait for 1000000 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8780 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 9460 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9000 ns;
channel_0 <= '0';
wait for 940 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8680 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9080 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 113870 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 8910 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 166090 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 9220 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 9320 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 61350 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 9160 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9270 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 61250 ns;
channel_0 <= '0';
wait for 960 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9050 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 61460 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61650 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8790 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 165930 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 61560 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 165480 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 140 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8780 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 420 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 26790 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 99470 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1600 ns;
channel_0 <= '1';
wait for 18260 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 90100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 570 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 1000000 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 311 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 599 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 501 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 9111 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 509 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 801 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 399 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 601 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 211 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 219 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 411 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 701 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 901 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 409 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 599 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 599 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9450 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 399 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 601 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 599 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 701 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 599 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 399 ns;
channel_0 <= '0';
wait for 401 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 939 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 401 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 701 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 389 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 119 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8581 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 120 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9089 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 389 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 309 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 409 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 489 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 311 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 113619 ns;
channel_0 <= '0';
wait for 731 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 491 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 191 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 309 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 909 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 89 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 89 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 409 ns;
channel_0 <= '0';
wait for 191 ns;
channel_0 <= '1';
wait for 8830 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 491 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 311 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 309 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 311 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 509 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 166110 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 911 ns;
channel_0 <= '1';
wait for 89 ns;
channel_0 <= '0';
wait for 911 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 909 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 399 ns;
channel_0 <= '1';
wait for 411 ns;
channel_0 <= '0';
wait for 589 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 399 ns;
channel_0 <= '1';
wait for 9291 ns;
channel_0 <= '0';
wait for 729 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 311 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 209 ns;
channel_0 <= '0';
wait for 191 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 499 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 699 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 601 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 309 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 309 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 601 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9340 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 389 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 309 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 911 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 909 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 389 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 701 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 610 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 389 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 409 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9249 ns;
channel_0 <= '0';
wait for 751 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 401 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 401 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 751 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 399 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 311 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 399 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 61250 ns;
channel_0 <= '0';
wait for 731 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 399 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 699 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 401 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 401 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 399 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 701 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 699 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9210 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 309 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 399 ns;
channel_0 <= '1';
wait for 211 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 191 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 191 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 401 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 911 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 509 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 491 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 909 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 909 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 399 ns;
channel_0 <= '1';
wait for 191 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 511 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 911 ns;
channel_0 <= '1';
wait for 89 ns;
channel_0 <= '0';
wait for 911 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 411 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 711 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 311 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 911 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 89 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 399 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 401 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 699 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9270 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 501 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 901 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 601 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 699 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 899 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 399 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 701 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 499 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 401 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 399 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 399 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 599 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 61199 ns;
channel_0 <= '0';
wait for 961 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 311 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 911 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 189 ns;
channel_0 <= '0';
wait for 610 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 411 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 399 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 191 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 191 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 9050 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 491 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 801 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 799 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 401 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 399 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 401 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 401 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 61480 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 401 ns;
channel_0 <= '1';
wait for 599 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 909 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 89 ns;
channel_0 <= '0';
wait for 311 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9249 ns;
channel_0 <= '0';
wait for 751 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 401 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 909 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 89 ns;
channel_0 <= '0';
wait for 911 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 401 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 609 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 899 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 901 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 9251 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 399 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 399 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 909 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 399 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 809 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 409 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 799 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 909 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 749 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 89 ns;
channel_0 <= '0';
wait for 111 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 909 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 311 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 811 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 499 ns;
channel_0 <= '0';
wait for 401 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 909 ns;
channel_0 <= '0';
wait for 191 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 191 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 111 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 399 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 701 ns;
channel_0 <= '1';
wait for 89 ns;
channel_0 <= '0';
wait for 111 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 399 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 89 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 749 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 89 ns;
channel_0 <= '0';
wait for 311 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 89 ns;
channel_0 <= '0';
wait for 311 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 909 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 311 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 89 ns;
channel_0 <= '0';
wait for 311 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 909 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 89 ns;
channel_0 <= '0';
wait for 911 ns;
channel_0 <= '1';
wait for 89 ns;
channel_0 <= '0';
wait for 911 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 909 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 909 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 89 ns;
channel_0 <= '0';
wait for 911 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 909 ns;
channel_0 <= '1';
wait for 91 ns;
channel_0 <= '0';
wait for 909 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61730 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 89 ns;
channel_0 <= '0';
wait for 911 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 309 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 8700 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 309 ns;
channel_0 <= '0';
wait for 81 ns;
channel_0 <= '1';
wait for 419 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 191 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 401 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 399 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 141 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 165619 ns;
channel_0 <= '0';
wait for 751 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 999 ns;
channel_0 <= '1';
wait for 61631 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 309 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 311 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 309 ns;
channel_0 <= '0';
wait for 491 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 309 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 899 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 309 ns;
channel_0 <= '0';
wait for 191 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 165399 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 901 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 191 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 409 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 211 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 309 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 149 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8780 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 409 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 311 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 391 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 201 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 889 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 891 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 189 ns;
channel_0 <= '1';
wait for 111 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 91 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 411 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 109 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 411 ns;
channel_0 <= '0';
wait for 89 ns;
channel_0 <= '1';
wait for 18521 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 301 ns;
channel_0 <= '0';
wait for 99 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 299 ns;
channel_0 <= '0';
wait for 301 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 599 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 799 ns;
channel_0 <= '1';
wait for 201 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 299 ns;
channel_0 <= '1';
wait for 401 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 99 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 199 ns;
channel_0 <= '0';
wait for 101 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 199 ns;
channel_0 <= '1';
wait for 101 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 108280 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1600 ns;
channel_0 <= '1';
wait for 117360 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1580 ns;
channel_0 <= '1';
wait for 225020 ns;
channel_0 <= '0';
wait for 960 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 3600 ns;
channel_0 <= '1';
wait for 1000000 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 140 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 9120 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 810 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9010 ns;
channel_0 <= '0';
wait for 940 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 710 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8680 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9090 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 113900 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 8880 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 165720 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9300 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9300 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 61330 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9220 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9270 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61200 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9040 ns;
channel_0 <= '0';
wait for 960 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 61480 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 490 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 390 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 710 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 710 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 9220 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61680 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 8780 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 165920 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 61620 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 165440 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9120 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9190 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 610 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9000 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 108440 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1600 ns;
channel_0 <= '1';
wait for 18250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 1000000 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9120 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 9100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9440 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9100 ns;
channel_0 <= '0';
wait for 940 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 610 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 810 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9080 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 113980 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 8800 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 166040 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9390 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9340 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 61210 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9270 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9270 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61150 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9040 ns;
channel_0 <= '0';
wait for 960 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 61460 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 9230 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61800 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 8670 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 320 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 165910 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 61700 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 165360 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 45100 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 7600 ns;
channel_0 <= '1';
wait for 63390 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 18340 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1600 ns;
channel_0 <= '1';
wait for 342000 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 3600 ns;
channel_0 <= '1';
wait for 1000000 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9440 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9000 ns;
channel_0 <= '0';
wait for 940 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 710 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 710 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 120 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8690 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9090 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 113880 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 8900 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 166030 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9300 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9330 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 61320 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9170 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9270 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 61240 ns;
channel_0 <= '0';
wait for 960 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9050 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 61460 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9230 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 990 ns;
channel_0 <= '1';
wait for 61710 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 8790 ns;
channel_0 <= '0';
wait for 880 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 165910 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61610 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 165450 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 120 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 570 ns;
channel_0 <= '1';
wait for 9560 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 108360 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1600 ns;
channel_0 <= '1';
wait for 18240 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 710 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 610 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 99480 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1580 ns;
channel_0 <= '1';
wait for 45030 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 3590 ns;
channel_0 <= '1';
wait for 1000000 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8780 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 140 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8780 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9430 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9090 ns;
channel_0 <= '0';
wait for 940 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 120 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 140 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8750 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 113960 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 8820 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 166020 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 290 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9390 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9340 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 61220 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9230 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 9240 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9270 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61190 ns;
channel_0 <= '0';
wait for 960 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9040 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 61460 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 760 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9230 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 61800 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 8690 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 165900 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61700 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 165380 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 580 ns;
channel_0 <= '1';
wait for 140 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 117220 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1590 ns;
channel_0 <= '1';
wait for 108370 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 6570 ns;
channel_0 <= '1';
wait for 9370 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 2600 ns;
channel_0 <= '1';
wait for 225020 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 3600 ns;
channel_0 <= '1';
wait for 1000000 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9470 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 8980 ns;
channel_0 <= '0';
wait for 940 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8690 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 9090 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 113880 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 8890 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 166030 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9300 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9300 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61360 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9190 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9240 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9280 ns;
channel_0 <= '0';
wait for 720 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 710 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 61240 ns;
channel_0 <= '0';
wait for 960 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9050 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61450 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1000 ns;
channel_0 <= '1';
wait for 61650 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 8790 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 165940 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61580 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 165450 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8770 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9380 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 117440 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1600 ns;
channel_0 <= '1';
wait for 18260 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 90100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 570 ns;
channel_0 <= '1';
wait for 140 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9230 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1600 ns;
channel_0 <= '1';
wait for 1000000 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 140 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8780 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9460 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9080 ns;
channel_0 <= '0';
wait for 940 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8600 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9090 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 113960 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 8810 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 166030 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9390 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9320 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 61260 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9230 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9270 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 61210 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9040 ns;
channel_0 <= '0';
wait for 960 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61440 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 610 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 61720 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 8710 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 165620 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61650 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 165380 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 140 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9320 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 610 ns;
channel_0 <= '1';
wait for 18270 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 18220 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 7600 ns;
channel_0 <= '1';
wait for 63360 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 18370 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1600 ns;
channel_0 <= '1';
wait for 107990 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 234270 ns;
channel_0 <= '0';
wait for 960 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 3600 ns;
channel_0 <= '1';
wait for 1000000 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 140 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9120 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 8980 ns;
channel_0 <= '0';
wait for 940 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 120 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8700 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 140 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8750 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8780 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 113890 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8880 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 166070 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9280 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9310 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61340 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 710 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9170 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9240 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 9270 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 710 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 61260 ns;
channel_0 <= '0';
wait for 960 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 9050 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61460 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9230 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61670 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 8790 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 80 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 165590 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 61610 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 165450 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 27130 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 99460 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1610 ns;
channel_0 <= '1';
wait for 18240 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 90120 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 570 ns;
channel_0 <= '1';
wait for 1000000 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 180 ns;
channel_0 <= '1';
wait for 8780 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9450 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9070 ns;
channel_0 <= '0';
wait for 940 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 8610 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 9080 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 113970 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 8810 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 150 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 165740 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9340 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9350 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9250 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 61220 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9210 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9240 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 800 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61200 ns;
channel_0 <= '0';
wait for 960 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 9040 ns;
channel_0 <= '0';
wait for 960 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 700 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 800 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61460 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 390 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 810 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 810 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 810 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 900 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 910 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 9260 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 410 ns;
channel_0 <= '1';
wait for 9220 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 61800 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 700 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 8670 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 510 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 165910 ns;
channel_0 <= '0';
wait for 750 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 61700 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 600 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 500 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 165370 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 610 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 790 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 690 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 9110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 390 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 18500 ns;
channel_0 <= '0';
wait for 740 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 110 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 490 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 190 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 610 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 210 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 810 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 600 ns;
channel_0 <= '1';
wait for 108310 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 190 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 210 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 310 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 710 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 710 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 910 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 410 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 510 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 310 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1600 ns;
channel_0 <= '1';
wait for 117370 ns;
channel_0 <= '0';
wait for 730 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 400 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 1580 ns;
channel_0 <= '1';
wait for 225030 ns;
channel_0 <= '0';
wait for 950 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 300 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 500 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 400 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 200 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 200 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 90 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 900 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 890 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 90 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 710 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 290 ns;
channel_0 <= '1';
wait for 110 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 590 ns;
channel_0 <= '1';
wait for 300 ns;
channel_0 <= '0';
wait for 100 ns;
channel_0 <= '1';
wait for 100 ns;
channel_0 <= '0';
wait for 3610 ns;
channel_0 <= '1';
    wait;
  end process;
end architecture;

